
   	